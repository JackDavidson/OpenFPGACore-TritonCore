module top(input a,input b, input c,input d, output x,output y);

assign x=a&b;
assign y=c&d;

endmodule
